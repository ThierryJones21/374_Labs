module control_unit(

output reg Gra,Grb, Grc, Rin, Rout, // here, you will define the inputs and outputs to your Control Unit
Yin, Zin,PCout, IncPC, MARin,Read, Write, Clear,ADD, AND, SHR,

input[31:0] IR, 
input Clock, Reset, Stop, Con_FF);           

parameter Reset_state= 4'b0000, fetch0 = 4'b0001, fetch1 = 4'b0010, fetch2= 4'b0011, add3 = 4'b0100, add4= 4'b0101, add5= 4'b0110;

reg [3:0] Present_state= Reset_state; // adjust the bit pattern based on the number of states

always@(posedge Clock, posedge Reset)// finite state machine; if clock or reset rising-edge
	begin if(Reset == 1'b1)
		Present_state =  Reset_state;
		else case(Present_state)
			Reset_state			:				Present_state = fetch0;
			
			fetch0				:				Present_state = fetch1;
			
			fetch1				:				Present_state = fetch2;
			fetch2				:				begin
														case(IR[31:27])   //inst. decoding based on the opcode to set the next state
															5'b00011:Present_state = add3;// this is the add instruction 
														endcase
													end
			add3					:				Present_state = add4;
			add4					:				Present_state = add5;
		endcase
	end
	
always@(Present_state)// do the job for each state
	begin case(Present_state)              // assert the required signals in each state
			Reset_state			:				begin Gra <= 0;   
														   Grb <= 0;  	 
															Grc <= 0; 
															Yin <= 0; //initialize the signals
													end
													
			fetch0				:				begin PCout<= 1; // see if you need to de-assert these signals 
															MARin <= 1;  
															IncPC <= 1; 
															Zin <= 0;
													end 
													
			add3					: 				begin Grb <= 1; 
															Rout<= 1;  
															Yin <= 0; 
													end
		endcase end
		
endmodule 