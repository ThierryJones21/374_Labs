module my374_lab1 ();
	reg temp;
endmodule 